library verilog;
use verilog.vl_types.all;
entity sync_fifo_tb is
end sync_fifo_tb;
