library verilog;
use verilog.vl_types.all;
entity async_fifo_tb is
end async_fifo_tb;
